/* until and s_until property */
/* property: as long as the RESET is high , CE should stay LOW */

module tb;
  
  reg clk = 0, rst = 0, ce = 0;
  always #5 clk = ~clk;
  
  
  initial begin
    rst = 1;
    #30;
    rst = 1;
    #10;
    ce = 0;
    rst = 1;
    #10;
    rst = 0;
    #50;
    ce = 0;
  end
  
  
  
  
  initial begin
    $dumpfile("dump.vcd"); 
    $dumpvars;
    $assertvacuousoff(0);
    #100;
    $finish();
  end
  
 initial A1: assert property (@(posedge clk) rst s_until ce) $info("Suc at %0t",$time);
 
endmodule
